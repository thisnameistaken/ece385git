module datapath();

endmodule