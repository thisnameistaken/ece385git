module top
(
    input   logic           Clk,        // 50MHz clock is only used to get timing estimate data
    input   logic           Reset,      // From push-button 0.  Remember the button is active low (0 when pressed)
    input   logic           ClearA_LoadB,      // From push-button 1
    input   logic           Run,        // From push-button 3.
    input   logic[7:0]      S,         // From slider switches
    
    // all outputs are registered
           
    output  logic[6:0]      AhexU,      
    output  logic[6:0]      AhexL,
    output  logic[6:0]      BhexU,
    output  logic[6:0]      BhexL,
    output  logic[7:0]      Aval,
    output  logic[7:0]      Bval,
	 output  logic           X
);

logic Reset_SH, ClrA_LdB, Run_SH;
logic [7:0] A, B, Din_S, sum;
logic x, add, sub, shift, clr_A, a_out, b_out, clr, cOut;

register_unit reg_unit(
							.Clk(Clk),
<<<<<<< HEAD
							.Reset(Reset_SH), //Button
							.X(x),
							.Add(add), 
							.Clr_Ld(clr),
							.Shift(shift),
							.ClearA(clr_A),
							.aout(a_out),
							.Ain(sum),
							.Bin(Din_S), //Switches
							.A_out(a_out),
							.B_out(b_out),
							.A(A),
							.B(B)
=======
							.Reset()
>>>>>>> 9eb7ff3ea75900aca39e99f23240c268b667bb17
							);

control c_unit(
				.Clk(Clk),
<<<<<<< HEAD
				.Reset(Reset_SH), //Button
				.Run(Run_SH), //Button
				.ClearA_LoadB(ClrA_LdB), 
				.x_in(x),
				.Bin(B),
				.Clr_Ld(clr),
				.Shift(shift),
				.Add(add),
				.Sub(sub),
				.X(x),
				.clearA(clr_A)
=======
				.Reset(),
				.Run(),
				.ClearA_LoadB(),
				.B(),
				.Clr_Ld(),
				.Shift(),
				.Add(),
				.Sub()
>>>>>>> 9eb7ff3ea75900aca39e99f23240c268b667bb17
				);

carry_select_adder adder_unit(
									.A(A),
									.B(Din_S),
									.A9(A[7]),
									.B9(Din_S[7]),
									.Sum(sum),
									.cOut(cOut),
									.X(x)
									);


HexDriver        HexAL (
                        .In0(A[3:0]),
                        .Out0(AhexL) );
HexDriver        HexBL (
                        .In0(B[3:0]),
                        .Out0(BhexL) );
HexDriver        HexAU (
                        .In0(A[6:3]),
                        .Out0(AhexU) );
HexDriver        HexBU (
                        .In0(B[6:3]),
                        .Out0(BhexU) );


	  //Input synchronizers required for asynchronous inputs (in this case, from the switches)
	  //These are array module instantiations
	  //Note: S stands for SYNCHRONIZED, H stands for active HIGH
	  //Note: We can invert the levels inside the port assignments
	  sync button_sync[3:0] (Clk, {~Reset, ~ClearA_LoadB, ~Run}, {Reset_SH, ClrA_LdB, Run_SH});
	  sync Din_sync[7:0] (Clk, Din, Din_S);

endmodule 